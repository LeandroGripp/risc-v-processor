LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

-- Instruction Memory, where it is stored the program in machine language
-- Built as a simple ROM memory
-- Instructions were translated from assembly code using riscV specifications
-- Instructions are stored during initialization, as we were not supposed to build a path for it to be stored

ENTITY InstructionMemory IS
  PORT (
    A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    RD : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END InstructionMemory;

ARCHITECTURE behavioral OF InstructionMemory IS
  TYPE ramType IS ARRAY(0 TO 26) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL ram : ramType := (--Initialize with assembly code translated into riscV machine code
  "00010000000000010000010100110111",
  "00001111100001010010010100000011",
  "00000000100000000000000011101111",
  "00000110000000000000000001101111",
  "00000000101000000000010000110011",
  "00000000001000000000001010010011",
  "00000010010101000110001100110011",
  "00000000000000110001101001100011",
  "00010000000000010000111000110111",
  "00001110010111100010111000100011",
  "00000010010101000100010000110011",
  "11111110110111111111000001101111",
  "00000000001100000000010010010011",
  "00000010100101001000001100110011",
  "00000010011001000100001001100011",
  "00000010100101000110001100110011",
  "00000000000000110001101001100011",
  "00010000000000010000111000110111",
  "00001110100111100010111000100011",
  "00000010100101000100010000110011",
  "11111110110111111111000001101111",
  "00000000010101001000010010110011",
  "11111101110111111111000001101111",
  "00000000010101000100011001100011",
  "00010000000000010000111000110111",
  "00001110100011100010111000100011",
  "00000000000000001000000001100111"
  );

  CONSTANT baseAddress : STD_LOGIC_VECTOR(31 DOWNTO 0) := x"00400000";

BEGIN
  PROCESS (A, ram) IS
    VARIABLE memIndex : INTEGER;
  BEGIN
    memIndex := to_integer((unsigned(A) - unsigned(baseAddress)) / 4);
    IF (memIndex <= 26) THEN
      RD <= ram(memIndex);
    ELSE
      RD <= x"00000000";
    END IF;
  END PROCESS;
END behavioral;